module VGA_Adjust_Speed(clk, rst, push, switch,	hsync, vsync, rgb);

input clk, rst;
input [1:0] push; 
input [2:0] switch;
output hsync, vsync;
output [2:0] rgb;

wire video_on;
wire [9:0] pixel_x, pixel_y;

// instantiate vgaSync and pixelGeneration circuit
//debounce debounce (.rst(rst), .clk(clk), .noisy(push), .clean(pushDB));
vgaSync vgaSync(.clk(clk), .rst(rst), .hsync(hsync), .vsync(vsync), .video_on(video_on), .p_tick(), .pixel_x(pixel_x), .pixel_y(pixel_y));

pixelGeneration pixelGeneration(.clk(clk), .rst(rst), .push(push), .switch(switch), .pixel_x(pixel_x), .pixel_y(pixel_y), .video_on(video_on), .rgb(rgb));

endmodule
